`define SIMULATION

module async_transmitter(
    input clk,
    input TxD_start,
    input [7:0] TxD_data,
    output TxD,
    output TxD_busy
);

// Assert TxD_start for (at least) one clock cycle to start transmission of TxD_data
// TxD_data is latched so that it doesn't have to stay valid while it is being sent
parameter ClkFrequency = 25000000; // 25MHz
parameter Baud = 115200;
parameter Oversampling = 1;        // Oversampling rate

`ifdef SIMULATION
    wire BitTick = 1'b1;  // output one bit per clock cycle
`else
    wire BitTick;

    BaudTickGen #(ClkFrequency, Baud, Oversampling) tickgen(
        .clk(clk),
        .enable(TxD_busy),
        .tick(BitTick)
    );
`endif

// Checks if frequency and baudate make sense
generate
    if (ClkFrequency < Baud * 8 && (ClkFrequency % Baud != 0)) ASSERTION_ERROR PARAMETER_OUT_OF_RANGE("Frequency incompatible with baud rate");
endgenerate


reg [3:0] TxD_state = 0;
reg [7:0] TxD_shift = 0;

wire TxD_ready = (TxD_state == 0);
assign TxD_busy = ~TxD_ready;

always @(posedge clk)
begin
    if(TxD_ready & TxD_start)
        TxD_shift <= TxD_data; // set TxD_shift to TxD_data
    else
        if(TxD_state[3] & BitTick)
            TxD_shift <= (TxD_shift >> 1); // shift right one bit

        case(TxD_state)
            4'b0000: if(TxD_start) TxD_state <= 4'b0100;
            4'b0100: if(BitTick) TxD_state <= 4'b1000;  // start bit
            4'b1000: if(BitTick) TxD_state <= 4'b1001;  // bit 0
            4'b1001: if(BitTick) TxD_state <= 4'b1010;  // bit 1
            4'b1010: if(BitTick) TxD_state <= 4'b1011;  // bit 2
            4'b1011: if(BitTick) TxD_state <= 4'b1100;  // bit 3
            4'b1100: if(BitTick) TxD_state <= 4'b1101;  // bit 4
            4'b1101: if(BitTick) TxD_state <= 4'b1110;  // bit 5
            4'b1110: if(BitTick) TxD_state <= 4'b1111;  // bit 6
            4'b1111: if(BitTick) TxD_state <= 4'b0010;  // bit 7
            4'b0010: if(BitTick) TxD_state <= 4'b0011;  // stop1
            4'b0011: if(BitTick) TxD_state <= 4'b0000;  // stop2
            default: if(BitTick) TxD_state <= 4'b0000;
        endcase
end

assign TxD = (TxD_state < 4) | (TxD_state[3] & TxD_shift[0]);  // put together the start, data and stop bits
endmodule
